class wzy_reg_reset_2_vseq extends uart_vseq_base;

`uvm_object_utils(wzy_reg_reset_2_vseq)

function new(string name = "wzy_reg_reset_vseq");
    super.new(name);
endfunction

task body;
    

endtask: body

endclass