module top_module( 
    input [3:0] in,
    output [2:0] out_both,
    output [3:1] out_any,
    output [3:0] out_different );
    
    integer i;
    
    always @(*) begin
        for(i = 0; i < 3; i ++) begin
            out_both[i] = in[i] & in[i+1];
            out_any[i+1] = in[i] | in[i+1];
            out_different[i] = (in[i] != in[i+1]) ? 1:0;
        end
        out_different[3] = (in[0] != in[3]) ? 1:0;
    end

endmodule
/*always @(*) begin
        for(int i = 0; i <= 3; i++) begin
            if(i <= 2)
                out_both[i] = in[i]&in[i+1];
            if(i >=1)
                out_any[i] = in[i]|in[i-1];
            
            if(i < 3)
                out_different[i] = in[i]^in[i+1];
            if(i ==3)
                out_different[3] = in[3]^in[0];
        end
    end
*/