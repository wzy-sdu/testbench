module soc_top (
    ports
);
    
endmodule