soc_top_clkrstn_intf()
logic m_sys_clk

`ifndef FPGA_EN
